library verilog;
use verilog.vl_types.all;
entity Relogio_tb is
end Relogio_tb;
